module SUM1BBC (A, B, Ci, Cout, S);

	input A;
	input B;
	input Ci;
	output Cout;
	output S;
	
	reg [1:0] st; //registro que guarda la suma
	assign S = st[0];
	assign Cout = st[1];
	//falta "<"
	always @ (*) begin
	st <= A+B+Ci;
	end 
	

endmodule

	